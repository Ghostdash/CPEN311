// nios_system_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_system_tb (
	);

	wire        nios_system_inst_clk_bfm_clk_clk;             // nios_system_inst_clk_bfm:clk -> [nios_system_inst:clk_clk, nios_system_inst_reset_bfm:clk]
	wire  [7:0] nios_system_inst_leds_export;                 // nios_system_inst:leds_export -> nios_system_inst_leds_bfm:sig_export
	wire  [7:0] nios_system_inst_switches_bfm_conduit_export; // nios_system_inst_switches_bfm:sig_export -> nios_system_inst:switches_export
	wire        nios_system_inst_reset_bfm_reset_reset;       // nios_system_inst_reset_bfm:reset -> nios_system_inst:reset_reset_n

	nios_system nios_system_inst (
		.clk_clk         (nios_system_inst_clk_bfm_clk_clk),             //      clk.clk
		.leds_export     (nios_system_inst_leds_export),                 //     leds.export
		.reset_reset_n   (nios_system_inst_reset_bfm_reset_reset),       //    reset.reset_n
		.switches_export (nios_system_inst_switches_bfm_conduit_export)  // switches.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nios_system_inst_clk_bfm (
		.clk (nios_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm nios_system_inst_leds_bfm (
		.sig_export (nios_system_inst_leds_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nios_system_inst_reset_bfm (
		.reset (nios_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nios_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 nios_system_inst_switches_bfm (
		.sig_export (nios_system_inst_switches_bfm_conduit_export)  // conduit.export
	);

endmodule
