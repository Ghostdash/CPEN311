// dnn_accel_system.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module dnn_accel_system (
		input  wire        clk_clk,           //        clk.clk
		output wire [6:0]  hex_export,        //        hex.export
		output wire        pll_locked_export, // pll_locked.export
		input  wire        reset_reset_n,     //      reset.reset_n
		output wire [12:0] sdram_addr,        //      sdram.addr
		output wire [1:0]  sdram_ba,          //           .ba
		output wire        sdram_cas_n,       //           .cas_n
		output wire        sdram_cke,         //           .cke
		output wire        sdram_cs_n,        //           .cs_n
		inout  wire [15:0] sdram_dq,          //           .dq
		output wire [1:0]  sdram_dqm,         //           .dqm
		output wire        sdram_ras_n,       //           .ras_n
		output wire        sdram_we_n,        //           .we_n
		output wire        sdram_clk_clk,     //  sdram_clk.clk
		output wire [7:0]  vga_vga_blu,       //        vga.vga_blu
		output wire        vga_vga_clk,       //           .vga_clk
		output wire [7:0]  vga_vga_grn,       //           .vga_grn
		output wire        vga_vga_hsync,     //           .vga_hsync
		output wire [7:0]  vga_vga_red,       //           .vga_red
		output wire        vga_vga_vsync      //           .vga_vsync
	);

	wire         pll_0_outclk0_clk;                                           // pll_0:outclk_0 -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_0_outclk0_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, pio_0:clk, rst_controller:clk, vga_avalon_0:clk, wordcopy_0:clk]
	wire  [31:0] wordcopy_0_avalon_master_readdata;                           // mm_interconnect_0:wordcopy_0_avalon_master_readdata -> wordcopy_0:master_readdata
	wire         wordcopy_0_avalon_master_waitrequest;                        // mm_interconnect_0:wordcopy_0_avalon_master_waitrequest -> wordcopy_0:master_waitrequest
	wire  [31:0] wordcopy_0_avalon_master_address;                            // wordcopy_0:master_address -> mm_interconnect_0:wordcopy_0_avalon_master_address
	wire         wordcopy_0_avalon_master_read;                               // wordcopy_0:master_read -> mm_interconnect_0:wordcopy_0_avalon_master_read
	wire         wordcopy_0_avalon_master_readdatavalid;                      // mm_interconnect_0:wordcopy_0_avalon_master_readdatavalid -> wordcopy_0:master_readdatavalid
	wire         wordcopy_0_avalon_master_write;                              // wordcopy_0:master_write -> mm_interconnect_0:wordcopy_0_avalon_master_write
	wire  [31:0] wordcopy_0_avalon_master_writedata;                          // wordcopy_0:master_writedata -> mm_interconnect_0:wordcopy_0_avalon_master_writedata
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [15:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;      // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;        // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;     // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;         // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;            // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;      // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;   // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;           // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;       // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_wordcopy_0_avalon_slave_readdata;          // wordcopy_0:slave_readdata -> mm_interconnect_0:wordcopy_0_avalon_slave_readdata
	wire         mm_interconnect_0_wordcopy_0_avalon_slave_waitrequest;       // wordcopy_0:slave_waitrequest -> mm_interconnect_0:wordcopy_0_avalon_slave_waitrequest
	wire   [3:0] mm_interconnect_0_wordcopy_0_avalon_slave_address;           // mm_interconnect_0:wordcopy_0_avalon_slave_address -> wordcopy_0:slave_address
	wire         mm_interconnect_0_wordcopy_0_avalon_slave_read;              // mm_interconnect_0:wordcopy_0_avalon_slave_read -> wordcopy_0:slave_read
	wire         mm_interconnect_0_wordcopy_0_avalon_slave_write;             // mm_interconnect_0:wordcopy_0_avalon_slave_write -> wordcopy_0:slave_write
	wire  [31:0] mm_interconnect_0_wordcopy_0_avalon_slave_writedata;         // mm_interconnect_0:wordcopy_0_avalon_slave_writedata -> wordcopy_0:slave_writedata
	wire  [31:0] mm_interconnect_0_vga_avalon_0_avalon_slave_0_readdata;      // vga_avalon_0:readdata -> mm_interconnect_0:vga_avalon_0_avalon_slave_0_readdata
	wire   [3:0] mm_interconnect_0_vga_avalon_0_avalon_slave_0_address;       // mm_interconnect_0:vga_avalon_0_avalon_slave_0_address -> vga_avalon_0:address
	wire         mm_interconnect_0_vga_avalon_0_avalon_slave_0_read;          // mm_interconnect_0:vga_avalon_0_avalon_slave_0_read -> vga_avalon_0:read
	wire         mm_interconnect_0_vga_avalon_0_avalon_slave_0_write;         // mm_interconnect_0:vga_avalon_0_avalon_slave_0_write -> vga_avalon_0:write
	wire  [31:0] mm_interconnect_0_vga_avalon_0_avalon_slave_0_writedata;     // mm_interconnect_0:vga_avalon_0_avalon_slave_0_writedata -> vga_avalon_0:writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;                       // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                         // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                          // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                            // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                        // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;            // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;              // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;               // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;            // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                 // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;             // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                 // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:wordcopy_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, onchip_memory2_0:reset, pio_0:reset_n, rst_translator:in_reset, vga_avalon_0:reset_n, wordcopy_0:rst_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	dnn_accel_system_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_0_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	dnn_accel_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (pll_0_outclk0_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                                //  wire.export
		.zs_ba          (sdram_ba),                                                  //      .export
		.zs_cas_n       (sdram_cas_n),                                               //      .export
		.zs_cke         (sdram_cke),                                                 //      .export
		.zs_cs_n        (sdram_cs_n),                                                //      .export
		.zs_dq          (sdram_dq),                                                  //      .export
		.zs_dqm         (sdram_dqm),                                                 //      .export
		.zs_ras_n       (sdram_ras_n),                                               //      .export
		.zs_we_n        (sdram_we_n)                                                 //      .export
	);

	dnn_accel_system_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_0_outclk0_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	dnn_accel_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_0_outclk0_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	dnn_accel_system_pio_0 pio_0 (
		.clk        (pll_0_outclk0_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (hex_export)                             // external_connection.export
	);

	dnn_accel_system_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.outclk_1 (sdram_clk_clk),     // outclk1.clk
		.locked   (pll_locked_export)  //  locked.export
	);

	vga_avalon vga_avalon_0 (
		.clk       (pll_0_outclk0_clk),                                       //          clock.clk
		.reset_n   (~rst_controller_reset_out_reset),                         //          reset.reset_n
		.address   (mm_interconnect_0_vga_avalon_0_avalon_slave_0_address),   // avalon_slave_0.address
		.read      (mm_interconnect_0_vga_avalon_0_avalon_slave_0_read),      //               .read
		.readdata  (mm_interconnect_0_vga_avalon_0_avalon_slave_0_readdata),  //               .readdata
		.write     (mm_interconnect_0_vga_avalon_0_avalon_slave_0_write),     //               .write
		.writedata (mm_interconnect_0_vga_avalon_0_avalon_slave_0_writedata), //               .writedata
		.vga_blu   (vga_vga_blu),                                             //    conduit_end.vga_blu
		.vga_clk   (vga_vga_clk),                                             //               .vga_clk
		.vga_grn   (vga_vga_grn),                                             //               .vga_grn
		.vga_hsync (vga_vga_hsync),                                           //               .vga_hsync
		.vga_red   (vga_vga_red),                                             //               .vga_red
		.vga_vsync (vga_vga_vsync)                                            //               .vga_vsync
	);

	wordcopy wordcopy_0 (
		.rst_n                (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.master_address       (wordcopy_0_avalon_master_address),                      // avalon_master.address
		.master_read          (wordcopy_0_avalon_master_read),                         //              .read
		.master_readdata      (wordcopy_0_avalon_master_readdata),                     //              .readdata
		.master_readdatavalid (wordcopy_0_avalon_master_readdatavalid),                //              .readdatavalid
		.master_waitrequest   (wordcopy_0_avalon_master_waitrequest),                  //              .waitrequest
		.master_write         (wordcopy_0_avalon_master_write),                        //              .write
		.master_writedata     (wordcopy_0_avalon_master_writedata),                    //              .writedata
		.slave_waitrequest    (mm_interconnect_0_wordcopy_0_avalon_slave_waitrequest), //  avalon_slave.waitrequest
		.slave_address        (mm_interconnect_0_wordcopy_0_avalon_slave_address),     //              .address
		.slave_read           (mm_interconnect_0_wordcopy_0_avalon_slave_read),        //              .read
		.slave_readdata       (mm_interconnect_0_wordcopy_0_avalon_slave_readdata),    //              .readdata
		.slave_write          (mm_interconnect_0_wordcopy_0_avalon_slave_write),       //              .write
		.slave_writedata      (mm_interconnect_0_wordcopy_0_avalon_slave_writedata),   //              .writedata
		.clk                  (pll_0_outclk0_clk)                                      //         clock.clk
	);

	dnn_accel_system_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                            (pll_0_outclk0_clk),                                           //                          pll_0_outclk0.clk
		.wordcopy_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // wordcopy_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address             (nios2_gen2_0_data_master_address),                            //               nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest         (nios2_gen2_0_data_master_waitrequest),                        //                                       .waitrequest
		.nios2_gen2_0_data_master_byteenable          (nios2_gen2_0_data_master_byteenable),                         //                                       .byteenable
		.nios2_gen2_0_data_master_read                (nios2_gen2_0_data_master_read),                               //                                       .read
		.nios2_gen2_0_data_master_readdata            (nios2_gen2_0_data_master_readdata),                           //                                       .readdata
		.nios2_gen2_0_data_master_write               (nios2_gen2_0_data_master_write),                              //                                       .write
		.nios2_gen2_0_data_master_writedata           (nios2_gen2_0_data_master_writedata),                          //                                       .writedata
		.nios2_gen2_0_data_master_debugaccess         (nios2_gen2_0_data_master_debugaccess),                        //                                       .debugaccess
		.nios2_gen2_0_instruction_master_address      (nios2_gen2_0_instruction_master_address),                     //        nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest  (nios2_gen2_0_instruction_master_waitrequest),                 //                                       .waitrequest
		.nios2_gen2_0_instruction_master_read         (nios2_gen2_0_instruction_master_read),                        //                                       .read
		.nios2_gen2_0_instruction_master_readdata     (nios2_gen2_0_instruction_master_readdata),                    //                                       .readdata
		.wordcopy_0_avalon_master_address             (wordcopy_0_avalon_master_address),                            //               wordcopy_0_avalon_master.address
		.wordcopy_0_avalon_master_waitrequest         (wordcopy_0_avalon_master_waitrequest),                        //                                       .waitrequest
		.wordcopy_0_avalon_master_read                (wordcopy_0_avalon_master_read),                               //                                       .read
		.wordcopy_0_avalon_master_readdata            (wordcopy_0_avalon_master_readdata),                           //                                       .readdata
		.wordcopy_0_avalon_master_readdatavalid       (wordcopy_0_avalon_master_readdatavalid),                      //                                       .readdatavalid
		.wordcopy_0_avalon_master_write               (wordcopy_0_avalon_master_write),                              //                                       .write
		.wordcopy_0_avalon_master_writedata           (wordcopy_0_avalon_master_writedata),                          //                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //          jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_0_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_0_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.new_sdram_controller_0_s1_address            (mm_interconnect_0_new_sdram_controller_0_s1_address),         //              new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write              (mm_interconnect_0_new_sdram_controller_0_s1_write),           //                                       .write
		.new_sdram_controller_0_s1_read               (mm_interconnect_0_new_sdram_controller_0_s1_read),            //                                       .read
		.new_sdram_controller_0_s1_readdata           (mm_interconnect_0_new_sdram_controller_0_s1_readdata),        //                                       .readdata
		.new_sdram_controller_0_s1_writedata          (mm_interconnect_0_new_sdram_controller_0_s1_writedata),       //                                       .writedata
		.new_sdram_controller_0_s1_byteenable         (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),      //                                       .byteenable
		.new_sdram_controller_0_s1_readdatavalid      (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),   //                                       .readdatavalid
		.new_sdram_controller_0_s1_waitrequest        (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),     //                                       .waitrequest
		.new_sdram_controller_0_s1_chipselect         (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),      //                                       .chipselect
		.nios2_gen2_0_debug_mem_slave_address         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //           nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                       .write
		.nios2_gen2_0_debug_mem_slave_read            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                       .read
		.nios2_gen2_0_debug_mem_slave_readdata        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                       .readdata
		.nios2_gen2_0_debug_mem_slave_writedata       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                       .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                       .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                       .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                       .debugaccess
		.onchip_memory2_0_s1_address                  (mm_interconnect_0_onchip_memory2_0_s1_address),               //                    onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                    (mm_interconnect_0_onchip_memory2_0_s1_write),                 //                                       .write
		.onchip_memory2_0_s1_readdata                 (mm_interconnect_0_onchip_memory2_0_s1_readdata),              //                                       .readdata
		.onchip_memory2_0_s1_writedata                (mm_interconnect_0_onchip_memory2_0_s1_writedata),             //                                       .writedata
		.onchip_memory2_0_s1_byteenable               (mm_interconnect_0_onchip_memory2_0_s1_byteenable),            //                                       .byteenable
		.onchip_memory2_0_s1_chipselect               (mm_interconnect_0_onchip_memory2_0_s1_chipselect),            //                                       .chipselect
		.onchip_memory2_0_s1_clken                    (mm_interconnect_0_onchip_memory2_0_s1_clken),                 //                                       .clken
		.pio_0_s1_address                             (mm_interconnect_0_pio_0_s1_address),                          //                               pio_0_s1.address
		.pio_0_s1_write                               (mm_interconnect_0_pio_0_s1_write),                            //                                       .write
		.pio_0_s1_readdata                            (mm_interconnect_0_pio_0_s1_readdata),                         //                                       .readdata
		.pio_0_s1_writedata                           (mm_interconnect_0_pio_0_s1_writedata),                        //                                       .writedata
		.pio_0_s1_chipselect                          (mm_interconnect_0_pio_0_s1_chipselect),                       //                                       .chipselect
		.vga_avalon_0_avalon_slave_0_address          (mm_interconnect_0_vga_avalon_0_avalon_slave_0_address),       //            vga_avalon_0_avalon_slave_0.address
		.vga_avalon_0_avalon_slave_0_write            (mm_interconnect_0_vga_avalon_0_avalon_slave_0_write),         //                                       .write
		.vga_avalon_0_avalon_slave_0_read             (mm_interconnect_0_vga_avalon_0_avalon_slave_0_read),          //                                       .read
		.vga_avalon_0_avalon_slave_0_readdata         (mm_interconnect_0_vga_avalon_0_avalon_slave_0_readdata),      //                                       .readdata
		.vga_avalon_0_avalon_slave_0_writedata        (mm_interconnect_0_vga_avalon_0_avalon_slave_0_writedata),     //                                       .writedata
		.wordcopy_0_avalon_slave_address              (mm_interconnect_0_wordcopy_0_avalon_slave_address),           //                wordcopy_0_avalon_slave.address
		.wordcopy_0_avalon_slave_write                (mm_interconnect_0_wordcopy_0_avalon_slave_write),             //                                       .write
		.wordcopy_0_avalon_slave_read                 (mm_interconnect_0_wordcopy_0_avalon_slave_read),              //                                       .read
		.wordcopy_0_avalon_slave_readdata             (mm_interconnect_0_wordcopy_0_avalon_slave_readdata),          //                                       .readdata
		.wordcopy_0_avalon_slave_writedata            (mm_interconnect_0_wordcopy_0_avalon_slave_writedata),         //                                       .writedata
		.wordcopy_0_avalon_slave_waitrequest          (mm_interconnect_0_wordcopy_0_avalon_slave_waitrequest)        //                                       .waitrequest
	);

	dnn_accel_system_irq_mapper irq_mapper (
		.clk           (pll_0_outclk0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
