// dnn_accel_system_tb.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module dnn_accel_system_tb (
	);

	wire         dnn_accel_system_inst_clk_bfm_clk_clk;             // dnn_accel_system_inst_clk_bfm:clk -> [dnn_accel_system_inst:clk_clk, dnn_accel_system_inst_reset_bfm:clk]
	wire         new_sdram_controller_0_my_partner_clk_bfm_clk_clk; // new_sdram_controller_0_my_partner_clk_bfm:clk -> new_sdram_controller_0_my_partner:clk
	wire   [6:0] dnn_accel_system_inst_hex_export;                  // dnn_accel_system_inst:hex_export -> dnn_accel_system_inst_hex_bfm:sig_export
	wire         dnn_accel_system_inst_pll_locked_export;           // dnn_accel_system_inst:pll_locked_export -> dnn_accel_system_inst_pll_locked_bfm:sig_export
	wire         dnn_accel_system_inst_sdram_cs_n;                  // dnn_accel_system_inst:sdram_cs_n -> new_sdram_controller_0_my_partner:zs_cs_n
	wire   [1:0] dnn_accel_system_inst_sdram_dqm;                   // dnn_accel_system_inst:sdram_dqm -> new_sdram_controller_0_my_partner:zs_dqm
	wire         dnn_accel_system_inst_sdram_cas_n;                 // dnn_accel_system_inst:sdram_cas_n -> new_sdram_controller_0_my_partner:zs_cas_n
	wire         dnn_accel_system_inst_sdram_ras_n;                 // dnn_accel_system_inst:sdram_ras_n -> new_sdram_controller_0_my_partner:zs_ras_n
	wire         dnn_accel_system_inst_sdram_we_n;                  // dnn_accel_system_inst:sdram_we_n -> new_sdram_controller_0_my_partner:zs_we_n
	wire  [12:0] dnn_accel_system_inst_sdram_addr;                  // dnn_accel_system_inst:sdram_addr -> new_sdram_controller_0_my_partner:zs_addr
	wire         dnn_accel_system_inst_sdram_cke;                   // dnn_accel_system_inst:sdram_cke -> new_sdram_controller_0_my_partner:zs_cke
	wire  [15:0] dnn_accel_system_inst_sdram_dq;                    // [] -> [dnn_accel_system_inst:sdram_dq, new_sdram_controller_0_my_partner:zs_dq]
	wire   [1:0] dnn_accel_system_inst_sdram_ba;                    // dnn_accel_system_inst:sdram_ba -> new_sdram_controller_0_my_partner:zs_ba
	wire   [7:0] dnn_accel_system_inst_vga_vga_grn;                 // dnn_accel_system_inst:vga_vga_grn -> dnn_accel_system_inst_vga_bfm:sig_vga_grn
	wire         dnn_accel_system_inst_vga_vga_vsync;               // dnn_accel_system_inst:vga_vga_vsync -> dnn_accel_system_inst_vga_bfm:sig_vga_vsync
	wire   [7:0] dnn_accel_system_inst_vga_vga_red;                 // dnn_accel_system_inst:vga_vga_red -> dnn_accel_system_inst_vga_bfm:sig_vga_red
	wire         dnn_accel_system_inst_vga_vga_clk;                 // dnn_accel_system_inst:vga_vga_clk -> dnn_accel_system_inst_vga_bfm:sig_vga_clk
	wire         dnn_accel_system_inst_vga_vga_hsync;               // dnn_accel_system_inst:vga_vga_hsync -> dnn_accel_system_inst_vga_bfm:sig_vga_hsync
	wire   [7:0] dnn_accel_system_inst_vga_vga_blu;                 // dnn_accel_system_inst:vga_vga_blu -> dnn_accel_system_inst_vga_bfm:sig_vga_blu
	wire         dnn_accel_system_inst_reset_bfm_reset_reset;       // dnn_accel_system_inst_reset_bfm:reset -> dnn_accel_system_inst:reset_reset_n

	dnn_accel_system dnn_accel_system_inst (
		.clk_clk           (dnn_accel_system_inst_clk_bfm_clk_clk),       //        clk.clk
		.hex_export        (dnn_accel_system_inst_hex_export),            //        hex.export
		.pll_locked_export (dnn_accel_system_inst_pll_locked_export),     // pll_locked.export
		.reset_reset_n     (dnn_accel_system_inst_reset_bfm_reset_reset), //      reset.reset_n
		.sdram_addr        (dnn_accel_system_inst_sdram_addr),            //      sdram.addr
		.sdram_ba          (dnn_accel_system_inst_sdram_ba),              //           .ba
		.sdram_cas_n       (dnn_accel_system_inst_sdram_cas_n),           //           .cas_n
		.sdram_cke         (dnn_accel_system_inst_sdram_cke),             //           .cke
		.sdram_cs_n        (dnn_accel_system_inst_sdram_cs_n),            //           .cs_n
		.sdram_dq          (dnn_accel_system_inst_sdram_dq),              //           .dq
		.sdram_dqm         (dnn_accel_system_inst_sdram_dqm),             //           .dqm
		.sdram_ras_n       (dnn_accel_system_inst_sdram_ras_n),           //           .ras_n
		.sdram_we_n        (dnn_accel_system_inst_sdram_we_n),            //           .we_n
		.sdram_clk_clk     (),                                            //  sdram_clk.clk
		.vga_vga_blu       (dnn_accel_system_inst_vga_vga_blu),           //        vga.vga_blu
		.vga_vga_clk       (dnn_accel_system_inst_vga_vga_clk),           //           .vga_clk
		.vga_vga_grn       (dnn_accel_system_inst_vga_vga_grn),           //           .vga_grn
		.vga_vga_hsync     (dnn_accel_system_inst_vga_vga_hsync),         //           .vga_hsync
		.vga_vga_red       (dnn_accel_system_inst_vga_vga_red),           //           .vga_red
		.vga_vga_vsync     (dnn_accel_system_inst_vga_vga_vsync)          //           .vga_vsync
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) dnn_accel_system_inst_clk_bfm (
		.clk (dnn_accel_system_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm dnn_accel_system_inst_hex_bfm (
		.sig_export (dnn_accel_system_inst_hex_export)  // conduit.export
	);

	altera_conduit_bfm_0002 dnn_accel_system_inst_pll_locked_bfm (
		.sig_export (dnn_accel_system_inst_pll_locked_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) dnn_accel_system_inst_reset_bfm (
		.reset (dnn_accel_system_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (dnn_accel_system_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0003 dnn_accel_system_inst_vga_bfm (
		.sig_vga_blu   (dnn_accel_system_inst_vga_vga_blu),   // conduit.vga_blu
		.sig_vga_clk   (dnn_accel_system_inst_vga_vga_clk),   //        .vga_clk
		.sig_vga_grn   (dnn_accel_system_inst_vga_vga_grn),   //        .vga_grn
		.sig_vga_hsync (dnn_accel_system_inst_vga_vga_hsync), //        .vga_hsync
		.sig_vga_red   (dnn_accel_system_inst_vga_vga_red),   //        .vga_red
		.sig_vga_vsync (dnn_accel_system_inst_vga_vga_vsync)  //        .vga_vsync
	);

	altera_sdram_partner_module new_sdram_controller_0_my_partner (
		.clk      (new_sdram_controller_0_my_partner_clk_bfm_clk_clk), //     clk.clk
		.zs_dq    (dnn_accel_system_inst_sdram_dq),                    // conduit.dq
		.zs_addr  (dnn_accel_system_inst_sdram_addr),                  //        .addr
		.zs_ba    (dnn_accel_system_inst_sdram_ba),                    //        .ba
		.zs_cas_n (dnn_accel_system_inst_sdram_cas_n),                 //        .cas_n
		.zs_cke   (dnn_accel_system_inst_sdram_cke),                   //        .cke
		.zs_cs_n  (dnn_accel_system_inst_sdram_cs_n),                  //        .cs_n
		.zs_dqm   (dnn_accel_system_inst_sdram_dqm),                   //        .dqm
		.zs_ras_n (dnn_accel_system_inst_sdram_ras_n),                 //        .ras_n
		.zs_we_n  (dnn_accel_system_inst_sdram_we_n)                   //        .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) new_sdram_controller_0_my_partner_clk_bfm (
		.clk (new_sdram_controller_0_my_partner_clk_bfm_clk_clk)  // clk.clk
	);

endmodule
